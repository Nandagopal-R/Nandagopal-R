`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 30.11.2022 16:06:46
// Design Name: 
// Module Name: pow
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module pow(clk);
wire [15:0] in;
reg [15:0] op;
reg [15:0] a[11:0],b[11:0],c[10:0],d,in1;
reg [15:0] y;
integer i,l;
input clk;


vio_0 in_out_name (
  .clk(clk),                // input wire clk
  .probe_in0(op),    // input wire [15 : 0] probe_in0
  .probe_out0(in)  // output wire [15 : 0] probe_out0
);

always @(posedge clk)
begin

a[0]=16'b00000000_00000000;   //0
a[1]=16'b00000000_00010000;  //0.0625
a[2]=16'b00000000_00011111;  //0.1211
a[3]=16'b00000000_00000000;   //0
a[4]=16'b00000000_00010000;  //0.0625
a[5]=16'b00000000_00011111;  //0.1211
a[6]=16'b00000000_00000000;   //0
a[7]=16'b00000000_00010000;  //0.0625
a[8]=16'b00000000_00011111;  //0.1211
a[9]=16'b00000000_00000000;   //0
a[10]=16'b00000000_00010000;  //0.0625
a[11]=16'b00000000_00011111;  //0.1211


b[0]=16'b00000000_00000000;  //0
b[1]=16'b00000100_00000000;  // 4 
b[2]=16'b00000011_00001011;  // 3.0457
b[3]=16'b00000000_00000000;  //0
b[4]=16'b00000100_00000000;  // 4 
b[5]=16'b00000011_00001011;  // 3.0457
b[6]=16'b00000000_00000000;  //0
b[7]=16'b00000100_00000000;  // 4 
b[8]=16'b00000011_00001011;  // 3.0457
b[9]=16'b00000000_00000000;  //0
b[10]=16'b00000100_00000000;  // 4 
b[11]=16'b00000011_00001011;  // 3.0457

c[0]=16'b01000000_00000000;  // 64
c[1]=16'b00010000_01001000;  //16.2849
c[2]=16'b01000000_00000000;  // 64
c[3]=16'b00010000_01001000;  //16.2849
c[4]=16'b01000000_00000000;  // 64
c[5]=16'b00010000_01001000;  //16.2849
c[6]=16'b01000000_00000000;  // 64
c[7]=16'b00010000_01001000;  //16.2849
c[8]=16'b01000000_00000000;  // 64
c[9]=16'b00010000_01001000;  //16.2849c[0]=16'b01000000_00000000;  // 64
c[10]=16'b00010000_01001000;  //16.2849

in1={8'b0,in[7:0]};

end

always @(posedge clk)
begin

if(in[15:8]==0)
d[15:0]=16'b00000001_0000000;
if(in[15:8]==1)
d[15:0]=16'b00000010_0000000;
if(in[15:8]==2)
d[15:0]=16'b00000100_0000000;
if(in[15:8]==3)
d[15:0]=16'b00001000_0000000;
if(in[15:8]==4)
d[15:0]=16'b00010000_0000000;
if(in[15:8]==5)
d[15:0]=16'b00100000_0000000;
if(in[15:8]==6)
d[15:0]=16'b01000000_0000000;
if(in[15:8]==2)
d[15:0]=16'b10000000_0000000;

for(i=0;i<=13;i=i+1)
begin
if(in1>=a[i] && in1<a[i+1])
l=i;
end

y=(b[l+1]-b[l])*(in1-a[l])/(a[l+1]-a[l])+b[l];
op=d*y;

end

endmodule
